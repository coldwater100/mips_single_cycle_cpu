`timescale 1ns/1ps

module tb_CP0();
    reg [31:0] Inst;
    reg [31:0] PCin;
    reg [31:0] Din;
    reg ExpSrc0, ExpSrc1, ExpSrc2;
    reg clk, enable, reset;
    wire ExRegWrite, IsEret, HasExp, ExpBlock;
    wire [31:0] PCout;
    wire [31:0] Dout;

    CP0 uut(
        .Inst(Inst),
        .PCin(PCin),
        .Din(Din),
        .ExpSrc0(ExpSrc0),
        .ExpSrc1(ExpSrc1),
        .ExpSrc2(ExpSrc2),
        .clk(clk),
        .enable(enable),
        .reset(reset),
        .ExRegWrite(ExRegWrite),
        .IsEret(IsEret),
        .HasExp(HasExp),
        .ExpBlock(ExpBlock),
        .PCout(PCout),
        .Dout(Dout)
    );

    // Clock generation
    initial clk = 0;
    always #5 clk = ~clk;

    task print_status;
    begin
        $display("Inst = 0x%08h", Inst);
        $display("PCin = 0x%08h", PCin);
        $display("Din  = 0x%08h", Din);
        $display("ExpSrc0 = %b, ExpSrc1 = %b, ExpSrc2 = %b", ExpSrc0, ExpSrc1, ExpSrc2);
        $display("ExRegWrite = %b", ExRegWrite);
        $display("IsEret     = %b", IsEret);
        $display("HasExp     = %b", HasExp);
        $display("ExpBlock   = %b", ExpBlock);
        $display("PCout      = 0x%08h", PCout);
        $display("Dout       = 0x%08h", Dout);
        $display("----------------------------------");
    end
    endtask

    task init;
    begin
        Inst = 32'h0;
        PCin = 32'h00400000;
        Din = 32'h12345678;
        ExpSrc0 = 0; ExpSrc1 = 0; ExpSrc2 = 0;
        enable = 0;
        reset = 1;
        #10; reset = 0;
        print_status();
    end
    endtask

    task exception_trigger_test;
    begin
        Inst = 32'h0;
        ExpSrc0 = 1;
        #10;
        ExpSrc0 = 0;
        #10;
        print_status();
    end
    endtask

    task epc_write_test;
    begin
        Inst = 32'h00000000; // sel=00, ExRegWrite=1
        ExpSrc0 = 0;
        enable = 0;
        #10;
        print_status();
    end
    endtask

    task epc_read_test;
    begin
        Inst = (2'b00 << 11); // sel = 00
        enable = 1;
        #10;
        print_status();
    end
    endtask

    task eret_test;
    begin
        Inst = 32'b010000_10000_00000_00000_00000_011000; // eret
        #10;
        print_status();
    end
    endtask

    initial begin
        $display("==== CP0 Module Testbench Start ====");

        $display("\n[Initialization]");
        init();

        $display("\n[Exception Trigger Test]");
        exception_trigger_test();

        $display("\n[EPC Write Test]");
        epc_write_test();

        $display("\n[EPC Read Test]");
        epc_read_test();

        $display("\n[ERET Instruction Test]");
        eret_test();

        #20;
        $display("==== CP0 Module Testbench Complete ====");
        $stop;
    end
endmodule

