
`timescale 1ns / 1ps

module tb_syscall_decoder;

    // ??
    reg clk;
    reg Enable;
    reg [31:0] v0;
    reg [31:0] a0;

    // ??
    wire Halt;
    wire [31:0] Hex;
    reg reset;

    // ??? ?? ????
    syscall_decoder uut (
        .clk(clk),
        .reset(reset),
        .Enable(Enable),
        .v0(v0),
        .a0(a0),
        .Halt(Halt),
        .Hex(Hex)
    );

    // ?? ??
    always #5 clk = ~clk;

    initial begin
        $display("--- Starting syscall_decoder Testbench ---");

        // ??? ??
	reset =1;
        clk = 0;
        Enable = 0;
        v0 = 0;
        a0 = 0;

        // Test 1: Enable = 1, v0 != 10 ? Halt = 0
        #10;
        Enable = 1;
        v0 = 32'd5;
        a0 = 32'h12345678;
        #10;
        $display("<Test 1: v0 != 10>");
        $display("v0 = 0x%08h, a0 = 0x%08h, Hex = 0x%08h, Halt = %b", v0, a0, Hex, Halt);

        // Test 2: Enable = 1, v0 == 10 ? Halt = 1
        v0 = 32'd10;  // syscall 10
        a0 = 32'hDEADBEEF;
        #10;
        $display("<Test 2: v0 == 10>");
        $display("v0 = 0x%08h, a0 = 0x%08h, Hex = 0x%08h, Halt = %b", v0, a0, Hex, Halt);

        // Test 3: Enable = 0 ? hex_reg ??, Halt = 0
        Enable = 0;
        v0 = 32'd10;
        a0 = 32'hAAAAAAAA;  // ? ?? ???? ??? ?
        #10;
        $display("<Test 3: Enable = 0>");
        $display("v0 = 0x%08h, a0 = 0x%08h, Hex = 0x%08h, Halt = %b", v0, a0, Hex, Halt);

        $display("--- End of Testbench ---");
        $stop;
    end

endmodule
