module tb_ctr_unit;
  reg [5:0] op, func;
  wire memread, memwrite, alusrc, jump, memtoreg, branch;
  wire regdst, regwrite, bneorbeq, isjal, zeroextend;
  wire readrs, readrt, issyscall, isjr, isshamt, iscop0;
  wire [3:0] aluop;

  ctr_unit dut(
    .op(op), .func(func),
    .memread(memread), .memwrite(memwrite), .alusrc(alusrc),
    .jump(jump), .memtoreg(memtoreg), .branch(branch),
    .regdst(regdst), .regwrite(regwrite), .bneorbeq(bneorbeq), .isjal(isjal), .zeroextend(zeroextend),
    .readrs(readrs), .readrt(readrt),
    .issyscall(issyscall), .isjr(isjr), .isshamt(isshamt), .iscop0(iscop0),
    .aluop(aluop)
  );

  initial begin
    $display("===== Control Unit Test Start =====");

    // LW
    op = 6'b100011; func = 6'bxxxxxx; #10;
    $display("LW (op=100011): memread=%b, alusrc=%b, memtoreg=%b, regwrite=%b", memread, alusrc, memtoreg, regwrite);

    // SW
    op = 6'b101011; func = 6'bxxxxxx; #10;
    $display("SW (op=101011): memwrite=%b, alusrc=%b", memwrite, alusrc);

    // R-type (ADD)
    op = 6'b000000; func = 6'b100000; #10;
    $display("R-type ADD (op=000000, func=100000): regdst=%b, regwrite=%b, aluop=%b", regdst, regwrite, aluop);

    // BEQ
    op = 6'b000100; func = 6'bxxxxxx; #10;
    $display("BEQ (op=000100): branch=%b, bneorbeq=%b", branch, bneorbeq);

    // BNE
    op = 6'b000101; func = 6'bxxxxxx; #10;
    $display("BNE (op=000101): branch=%b, bneorbeq=%b", branch, bneorbeq);

    // JAL
    op = 6'b000011; func = 6'bxxxxxx; #10;
    $display("JAL (op=000011): jump=%b, isjal=%b, regwrite=%b", jump, isjal, regwrite);

    // LUI
    op = 6'b001111; func = 6'bxxxxxx; #10;
    $display("LUI (op=001111): zeroextend=%b", zeroextend);

    // SYSCALL
    op = 6'b000000; func = 6'b001100; #10;
    $display("SYSCALL (op=000000, func=001100): issyscall=%b", issyscall);

    // JR
    op = 6'b000000; func = 6'b001000; #10;
    $display("JR (op=000000, func=001000): isjr=%b", isjr);

    // SLL
    op = 6'b000000; func = 6'b000000; #10;
    $display("SLL (op=000000, func=000000): isshamt=%b", isshamt);

    // COP0
    op = 6'b010000; func = 6'bxxxxxx; #10;
    $display("COP0 (op=010000): iscop0=%b", iscop0);

    $display("===== Control Unit Test End =====");
    $stop;
  end
endmodule

