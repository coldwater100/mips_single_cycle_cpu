`timescale 1ns / 1ps

module tb_instruction_memory;

    // ??
    reg [31:0] pc;

    // ??
    wire [31:0] data;

    // ??? ?? ?? ?????
    instruction_memory uut (
        .pc(pc),
        .data(data)
    );

    initial begin
        $display("\n=== Instruction Memory Testbench ===\n");

        // ???
        pc = 32'h00000000;
        #10 $display("pc = 0x%08h, data = 0x%08h", pc, data);

        pc = 32'h00000004;
        #10 $display("pc = 0x%08h, data = 0x%08h", pc, data);

        pc = 32'h00000008;
        #10 $display("pc = 0x%08h, data = 0x%08h", pc, data);

        pc = 32'h00000800; // sel = 1, rom1?? ?? ??
        #10 $display("pc = 0x%08h, data = 0x%08h", pc, data);

        pc = 32'h00000804;
        #10 $display("pc = 0x%08h, data = 0x%08h", pc, data);

        pc = 32'h00000808;
        #10 $display("pc = 0x%08h, data = 0x%08h", pc, data);

        $display("\n=== Testbench End ===");
        $stop;
    end

endmodule

