module mux #(
    // ?? ?? ? (? ?? ?? ? ???? ??)
    parameter integer select_bit = 2,
    // ? ?? ???? ?
    parameter integer data_bits   = 8
)(
    input  wire [select_bit-1:0]                     sel,       // ?? ??
    input  wire [(1<<select_bit)*data_bits-1:0]      data_bus,  // 2^select_bit?? data_bits ? ??? ??? ??? ??
    output reg  [data_bits-1:0]                      out        // ??? ??? ????
);

    integer i;
    always @* begin
        // ??? (0) ??
        out = {data_bits{1'b0}};
        // ?? ?? ??? ???? sel ?? ???? ???? ????? ??
        for (i = 0; i < (1<<select_bit); i = i + 1) begin
            if (sel == i) begin
                // SystemVerilog ??? ?? ?????: [base +: width]
                out = data_bus[i*data_bits +: data_bits];
            end
        end
    end

endmodule

